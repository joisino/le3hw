module core( input logic         clk,
            input logic         reset,

            input logic [15:0]  in_dat,
            output logic        out_en,
            output logic [15:0] out_dat,
            output logic        is_halt,

            output logic [15:0] pc,
            input logic [15:0]  inst,

            output logic [15:0] main_mem_read_adr,
            input logic [15:0]  main_mem_dat,
            output logic        main_mem_write,
            output logic [15:0] main_mem_write_adr,
            output logic [15:0] main_mem_write_dat );

   logic [15:0] pcinc, pcinc_id, pcinc_ex;
   logic [15:0] inst_id;
   logic [15:0] rd1_id, rd1_ex, rd1_mem, rd1_wb;
   logic [15:0] rd2_id, rd2_ex;
   logic [3:0]  d_id, d_ex;
   logic [15:0] extended_d_id, extended_d_ex, extended_d_mem, extended_d_wb;
   logic [2:0]  regwrite_adr_id, regwrite_adr_ex, regwrite_adr_mem;
   logic [1:0]  ALUsrcA_controll_id, ALUsrcA_controll;
   logic [1:0]  ALUsrcB_controll_id, ALUsrcB_controll;
   logic [3:0]  ALUop_id, ALUop;
   logic        main_mem_write_id, main_mem_write_ex;
   logic        regwrite_id, regwrite_ex, regwrite_mem, regwrite;
   logic        regwrite_dat_controll_id, regwrite_dat_controll_ex, regwrite_dat_controll_mem, regwrite_dat_controll;
   logic [15:0] ALUres_ex, ALUres_mem, ALUres_wb;
   logic        S_ex, S_mem, S_wb;
   logic        C_ex, C_mem, C_wb;
   logic        Z_ex, Z_mem, Z_wb;
   logic        V_ex, V_mem, V_wb;
   
   fetch fetch( .* );
   
   ifid ifid( .* );

   decode decode( .* );

   idex idex( .* );

   exec exec( .* );

   exmem exmem( .* );

   mainmem mainmem( .* );

   memwb memwb( .* );

   writeback writeback( .* );
   
endmodule
   
